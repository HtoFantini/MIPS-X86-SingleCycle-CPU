-- PORTA AND

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

-- RAM entity
ENTITY PORTA_AND IS
PORT(
       INPUT_1 : IN STD_LOGIC;
       INPUT_2 : IN STD_LOGIC;
       OUTPUT: OUT STD_LOGIC
    );
END ENTITY;

-- RAM architecture
ARCHITECTURE BEV OF PORTA_AND IS
BEGIN

	OUTPUT <= INPUT_1 AND INPUT_2;
    
END BEV;

