-- ALU CONTROL

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

-- ALU CONTROL ENTITY
ENTITY ALU_CONTROL IS
    PORT(
       ALU_OP : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
       BIT_30 : IN STD_LOGIC;
       BIT_14_12 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
       OPERATION : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END ENTITY;


ARCHITECTURE BEV OF ALU_CONTROL IS
BEGIN
	PROCESS(ALU_OP, BIT_30, BIT_14_12)
    BEGIN
	 
	 
		IF(ALU_OP = "011") THEN
			IF(BIT_14_12 = "000") THEN		--BEQ
				OPERATION <= "1111";
				ELSIF(BIT_14_12 = "101") THEN	--BGE
				OPERATION <= "0111";
				END IF;	--COMPLETAR COM OUTRAS INSTRUÇÕES DE BRANCH (TIPO B)
			
		ELSIF(ALU_OP = "101") THEN			--JALR
			OPERATION <= "1101";
		
		ELSIF(ALU_OP = "100") THEN			--TIPO I
			IF(BIT_14_12 = "000") THEN	    --ADDI
				OPERATION <="0010";
			ELSIF (BIT_14_12 = "001") THEN	--SLLI
				OPERATION <="0010";
			ELSIF (BIT_14_12 = "010") THEN	--SLTI
				OPERATION <="0010";
			ELSIF (BIT_14_12 = "011") THEN	--SLTIU
				OPERATION <="0010";
			ELSIF (BIT_14_12 = "100") THEN	--XORI
				OPERATION <="0010";
			ELSIF (BIT_14_12 = "101") THEN
				IF(BIT_30 = '0') THEN		--SRLI
					OPERATION <= "0011";
				ELSE						--SRAI
					OPERATION <="0010";
				END IF;
			ELSIF (BIT_14_12 = "110") THEN	--ORI
				OPERATION <="0001";
			ELSIF (BIT_14_12 = "111") THEN	--ANDI
				OPERATION <="0000";
			ELSE
				OPERATION <= "1111";
			END IF;
		ELSE
			IF (ALU_OP = "000") THEN
				 OPERATION <= "0010";
			ELSIF (ALU_OP(0) = '1') THEN
				 OPERATION <= "0110";
			ELSIF ((ALU_OP(1) = '1') AND (BIT_30 = '0') AND (BIT_14_12 = "000")) THEN
				 OPERATION <= "0010";
			ELSIF ((ALU_OP(1) = '1') AND (BIT_30 = '1') AND (BIT_14_12 = "000")) THEN
				 OPERATION <= "0010";
			ELSIF ((ALU_OP(1) = '1') AND (BIT_30 = '0') AND (BIT_14_12 = "111")) THEN
				 OPERATION <= "0000";
			ELSIF ((ALU_OP(1) = '1') AND (BIT_30 = '0') AND (BIT_14_12 = "110")) THEN
				 OPERATION <= "0001";
			ELSE
				 OPERATION <= "ZZZZ";
			END IF;
					
		END IF;

    
    END PROCESS;
END BEV;





